localparam A1_ADDRWIDTH = 9;
localparam A1_DATAWIDTH = 18;
localparam B1_ADDRWIDTH = A1_ADDRWIDTH;
localparam B1_DATAWIDTH = A1_DATAWIDTH;


localparam A2_ADDRWIDTH = 9;
localparam A2_DATAWIDTH = 18;
localparam B2_ADDRWIDTH = A2_ADDRWIDTH;
localparam B2_DATAWIDTH = A2_DATAWIDTH;

localparam DEPTH1 = 2**A1_ADDRWIDTH;
localparam DEPTH2 = 2**A1_ADDRWIDTH;

localparam BYTEWIDTH = 9;