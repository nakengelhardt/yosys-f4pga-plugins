localparam ABITS_A = 10;
localparam DBITS_A = 36;

localparam ABITS_B = ABITS_A;
localparam DBITS_B = DBITS_A;

localparam DEPTH = 2**(ABITS_A);
