localparam ABITS = 8;
localparam DBITS = 32;

localparam DEPTH = 2**ABITS;

localparam BYTEWIDTH = 8;
localparam NBYTES = DBITS/BYTEWIDTH;
