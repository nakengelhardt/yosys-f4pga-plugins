localparam ABITS = 10;
localparam DBITS = 18;

localparam DEPTH = 2**(ABITS+1);
