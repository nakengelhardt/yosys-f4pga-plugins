localparam ABITS = 10;
localparam DBITS = 18;

localparam DEPTH = 2**ABITS;

localparam BYTEWIDTH = 9;
localparam NBYTES = DBITS/BYTEWIDTH;