localparam ABITS = 12;
localparam DBITS = 8;

localparam DEPTH = 2**ABITS;
