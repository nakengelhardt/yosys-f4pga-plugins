localparam WABITS = 12;
localparam WDBITS = 9;

localparam RABITS = WABITS;
localparam RDBITS = WDBITS;

localparam DEPTH = 2**(WABITS+1);
