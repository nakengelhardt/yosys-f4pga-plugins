localparam ABITS = 9;
localparam DBITS = 18;

localparam DEPTH = 2**(ABITS+1);

localparam BYTEWIDTH = 9;
localparam NBYTES = DBITS/BYTEWIDTH;
